   // SSD
   output [3:0] ssd_anode,
   output       ssd_dp,		
   output [6:0] ssd_seg,
		
		
