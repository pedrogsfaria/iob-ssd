/*
 * file    hex2ssd.v
 * date    December 2022
 * 
 * brief   Seven-Segment Display (SSD) decoder.
 *         Converts a binary-coded decimal (BCD) to 7-bits SSD.  
*/
`timescale 1ns/1ps

module hex2ssd  
   (
    input [3:0]      bcd_number,    
    output reg [6:0] seg 
    );

   always @(*)
     begin
	case (bcd_number)
	  4'b0000: seg = 7'b1111110; // 0 
	  4'b0001: seg = 7'b0110000; // 1 
	  4'b0010: seg = 7'b1101101; // 2 
	  4'b0011: seg = 7'b1111001; // 3
	  4'b0100: seg = 7'b0110011; // 4 
          4'b0101: seg = 7'b0100100; // 5 
          4'b0110: seg = 7'b0100000; // 6 
          4'b0111: seg = 7'b0001111; // 7
          4'b1000: seg = 7'b0000000; // 8     
          4'b1001: seg = 7'b0000100; // 9    
	  4'b1010: seg = 7'b0000010; // A
	  4'b1011: seg = 7'b1100000; // B
	  4'b1100: seg = 7'b0110001; // C
	  4'b1101: seg = 7'b1000010; // D
	  4'b1110: seg = 7'b0110000; // E
	  4'b1111: seg = 7'b0111000; // F
          default: seg = 7'b0000001; // 0: 4b'0000
	endcase // case (bcd_number)
     end // always @ (*)

endmodule // hex2ssd
