   // SSD
   // input [13:0] ssd_data_in,
   output [3:0] ssd_anode,
   output [7:0] ssd_seg,
